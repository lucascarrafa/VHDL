LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY Decoder IS PORT(
	E: IN STD_LOGIC; 
	A: IN STD_LOGIC_VECTOR(2 DOWNTO 0); 
	Y: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)); 
END Decoder;
ARCHITECTURE Behavioral OF Decoder IS
BEGIN
 PROCESS (E, A)
 BEGIN
	 IF (E = '0') THEN 
		Y <= (OTHERS => '0'); 
	 ELSE
		 CASE A IS 
			 WHEN "000" => Y <= "00000001";
			 WHEN "001" => Y <= "00000010";
			 WHEN "010" => Y <= "00000100";
			 WHEN "011" => Y <= "00001000";
			 WHEN "100" => Y <= "00010000";
			 WHEN "101" => Y <= "00100000";
			 WHEN "110" => Y <= "01000000";
			 WHEN "111" => Y <= "10000000";
			 WHEN OTHERS => NULL;
		 END CASE;
	 END IF;
 END PROCESS;
END Behavioral; 